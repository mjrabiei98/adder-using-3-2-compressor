LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY adder6tw2 IS
    GENERIC (BITS : INTEGER := 8);
    PORT (
        op1, op2, op3, op4, op5, op6 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        OUT0 : OUT STD_LOGIC_VECTOR (BITS + 1 DOWNTO 0);
        OUT1 : OUT STD_LOGIC_VECTOR (BITS + 1 DOWNTO 0)
    );
END ENTITY;


ARCHITECTURE linear OF adder6tw2 IS
    SIGNAL w1 : STD_LOGIC_VECTOR(BITS - 1 DOWNTO 0);
    SIGNAL w2 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w3 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w4 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL w5 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w6 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL w7 : STD_LOGIC_VECTOR(BITS + 2 DOWNTO 0);
    SIGNAL t1 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL t2 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL t3 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL t4 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL t5 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
BEGIN
    t1 <= ('0' & op3);
    t2 <= ('0' & w1);
    t3 <= ('0' & op2);
    t4 <= ("00" & op1);
    t5 <= ('0' & w5);
    UI1 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS) PORT MAP(op6, op5, op4, w1, w2);
    UI2 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS + 1) PORT MAP(t1, t2, w2, w3, w4);
    UI3 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS + 1) PORT MAP(t3, w3, w4(BITS DOWNTO 0), w5, w6);
    UI4 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS + 2) PORT MAP(t4, t5, w6, OUT0, w7);
    OUT1 <= w7(BITS + 1 DOWNTO 0);
END ARCHITECTURE;

--------------------------------

ARCHITECTURE adder_tree OF adder6tw2 IS
    SIGNAL w1 : STD_LOGIC_VECTOR(BITS - 1 DOWNTO 0);
    SIGNAL w2 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w3 : STD_LOGIC_VECTOR(BITS - 1 DOWNTO 0);
    SIGNAL w4 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w5 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL w6 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL w7 : STD_LOGIC_VECTOR(BITS + 2 DOWNTO 0);
    SIGNAL t1 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
    SIGNAL t2 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL t3 : STD_LOGIC_VECTOR(BITS + 1 DOWNTO 0);
    SIGNAL t4 : STD_LOGIC_VECTOR(BITS DOWNTO 0);
BEGIN
    t1 <= ('0' & w3);
    t2 <= ('0' & w4);
    t3 <= ('0' & w5);
    t4 <= ('0' & w1);
    UI1 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS) PORT MAP(op6, op5, op4, w1, w2);
    UI2 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS) PORT MAP(op3, op2, op1, w3, w4);
    UI3 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS + 1) PORT MAP(t1, t4, w2, w5, w6);
    UI4 : ENTITY WORK.compressor3_2 GENERIC MAP(BITS + 2) PORT MAP(t2, t3, w6, OUT0, w7);
    OUT1 <= w7(BITS + 1 DOWNTO 0);
END ARCHITECTURE;